../../adder.vhd